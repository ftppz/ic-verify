// alu_pkg.sv

package alu_pkg;

  import rpt_pkg::*;

  `include "trans.sv"

  `include "generator.sv"

  `include "driver.sv"

  `include "monitor.sv"

  `include "agent.sv"
  
  `include "refmod.sv"

  `include "checker.sv"

  `include "coverage.sv"

  `include "env.sv"
  
  `include "base_test.sv"
  
  
endpackage:alu_pkg
